** Profile: "SCHEMATIC1-pr42"  [ C:\PROGRAM FILES\ORCAD\CAPTURE\PROJECTS\SCHEMATA4\pr4-SCHEMATIC1-pr42.sim ] 

** Creating circuit file "pr4-SCHEMATIC1-pr42.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN TEMP -20 130 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pr4-SCHEMATIC1.net" 


.END
