** Profile: "SCHEMATIC1-pr3"  [ c:\PROGRAM FILES\ORCAD\CAPTURE\PROJECTS\schemata3-SCHEMATIC1-pr3.sim ] 

** Creating circuit file "schemata3-SCHEMATIC1-pr3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\schemata3-SCHEMATIC1.net" 


.END
