** Profile: "SCHEMATIC1-pr12"  [ D:\�������\����������\������������\DSK\Prz\Orcad pr\SCHEMATA1\pr1-schematic1-pr12.sim ] 

** Creating circuit file "pr1-schematic1-pr12.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN TEMP -20 70 1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pr1-SCHEMATIC1.net" 


.END
