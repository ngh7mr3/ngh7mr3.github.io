** Profile: "SCHEMATIC1-pr21"  [ C:\PROGRAM FILES\ORCAD\CAPTURE\PROJECTS\SCHEMATA2\pr2-SCHEMATIC1-pr21.sim ] 

** Creating circuit file "pr2-SCHEMATIC1-pr21.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pr2-SCHEMATIC1.net" 


.END
