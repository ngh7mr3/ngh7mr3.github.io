** Profile: "SCHEMATIC1-pr43"  [ C:\PROGRAM FILES\ORCAD\CAPTURE\PROJECTS\SCHEMATA4\pr4-SCHEMATIC1-pr43.sim ] 

** Creating circuit file "pr4-SCHEMATIC1-pr43.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pr4-SCHEMATIC1.net" 


.END
